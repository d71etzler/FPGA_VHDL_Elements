--------------------------------------------------------------------------------
-- File: tb_func_spi.vhd
--
-- !THIS FILE IS UNDER REVISION CONTROL!
--
-- $Author:: uid03580  $: Author of last commit
-- $Date:: 2017-03-01 #$: Date of last commit
-- $Rev:: 34           $: Revision of last commit
--
-- Open Points/Remarks:
--  + (none)
--
--------------------------------------------------------------------------------

--------------------------------------------------------------------------------
-- Used library definitions
--------------------------------------------------------------------------------
library ieee;
  use ieee.numeric_std.all;
  use ieee.std_logic_1164.all;
  use ieee.std_logic_textio.all;
library spi;
  use spi.spi_elements.all;
library std;
  use std.textio.all;

--------------------------------------------------------------------------------
-- Package declarations
--------------------------------------------------------------------------------
package tb_func_spi is

--------------------------------------------------------------------------------
-- User constants
--------------------------------------------------------------------------------
-- (none)

--------------------------------------------------------------------------------
-- Type declarations
--------------------------------------------------------------------------------
-- (none)

--------------------------------------------------------------------------------
-- Function declarations
--------------------------------------------------------------------------------
-- (none)

end package tb_func_spi;

--------------------------------------------------------------------------------
-- Package definitions
--------------------------------------------------------------------------------
package body tb_func_spi is
end package body tb_func_spi;
